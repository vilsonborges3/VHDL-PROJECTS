
--PRODETO DE UM CIRCUITO LOGICO COMBNACIONAL 

ENTITY CIRCUITO1 IS
PORT (A, B, C, D : IN BIT;
	  S          : OUT BIT );
END CIRCUITO1;

ARCHITECTURE CIR OF CIRCUITO1 IS
BEGIN

S <=(( NOT ( A AND B AND C )) OR ( NOT C )) XOR ( C AND D ) ;
END CIR;