
--PROJETO DMUX 1X4

ENTITY M12011EAU020 IS
PORT (D, A, B : IN BIT ;
		S0, S1, S2, S3: OUT BIT );
END M12011EAU020 ;

ARCHITECTURE CIR OF M12011EAU020 IS 
SIGNAL VAR : BIT_VECTOR (1 DOWNTO 0) ;

BEGIN 
VAR <= A & B;

S0 <= D WHEN VAR = "00" ELSE '0';
S1 <= D WHEN VAR = "01" ELSE '0';
S2 <= D WHEN VAR = "10" ELSE '0';
S3 <= D WHEN VAR = "11" ELSE '0';

END CIR;