-- IMPLEMENTACAO DE UMA PORTA LOGICA E UTILIZANDO VHDL 

ENTITY PORTAS1 IS

PORT (A, B: IN BIT;
		S: OUT BIT);
		
END PORTAS1;

ARCHITECTURE CIRC OF PORTAS1 IS
BEGIN
 S <= A AND B ;
 END CIRC; 
