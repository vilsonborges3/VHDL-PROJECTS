--PROJETO FLIPFLOPJK MESTRE-ESCRAVO

ENTITY FLIPFLOP IS
PORT (PRN, CLRN, CLKN, J, K : IN BIT;
	Q : BUFFER BIT );
END FLIPFLOP;

ARCHITECTURE CIR OF FLIPFLOP IS

BEGIN

	PROCESS( PRN, CLRN, CLKN )
	BEGIN 
		IF PRN = '0' THEN Q <= '1';
		ELSIF CLRN = '0' THEN Q <= '0';
		ELSIF CLKN = '0' AND CLKN 'EVENT THEN 
			IF J = '1' AND K = '1' THEN Q <= NOT Q;
			ELSIF J = '1' AND K = '0' THEN Q <= '1';
			ELSIF J = '0' AND K = '1' THEN Q <= '0';
			END IF;
		END IF;
	END PROCESS;
	Q<=Q;
END CIR;
		
			
			
		
		
		
		
--CLK = BAIXO, ALTO, BORDA DE DESCIDA , BORDA DE SUBIDA 

--IF CLK='0' THEN (NIVEL BAIXO)
--IF CLK='1' THEN (NIVEL ALTO)
--PRA TESTAR BRDA USA EVENTO DE DECIDA OU SUBIDA:
--IF CLK = '0' AND CLK 'EVENT 