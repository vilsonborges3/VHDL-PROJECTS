ENTITY TRABALHO02 IS
PORT (A, B, C, D : IN BIT;
      S          : OUT BIT);
END TRABALHO02;

ARCHITECTURE CIR OF TRABALHO02 IS 
BEGIN 

S <= NOT( ( NOT( NOT( A AND (NOT C) AND D) OR ((NOT A) OR B OR (NOT C)) ) AND ( NOT C )) OR (B XOR D) OR ( NOT(((NOT A) OR B OR (NOT C)) AND D)) );
END CIR;