ENTITY M12011EAU020 IS 
PORT (A, B, C, D : IN BIT ;
      S          : OUT BIT );
END M12011EAU020 ;

ARCHITECTURE CIR OF M12011EAU020 IS 

SIGNAL S1, S2, S3, S4, S5, S6 : BIT;

BEGIN 

S <= NOT (S1 OR S6 OR S5);

S6 <= S4 AND (NOT C) ;
S5 <= NOT ((NOT S3) AND D) ;
S4 <= NOT (S2 OR S3) ;
S1 <= B XOR D;
S2 <= NOT(A AND (NOT C) AND D) ;
S3 <= NOT ((NOT A) OR B OR (NOT C));

END CIR;