-- PROJETO DE UM MUX 4X1

ENTITY M12011EAU020 IS
PORT ( D : IN BIT_VECTOR (3 DOWNTO 0) ;
       VAR : INTEGER RANGE 0 TO 3;
       S : OUT BIT);
END M12011EAU020 ;

ARCHITECTURE CIR OF M12011EAU020 IS 

BEGIN 

WITH VAR SELECT 

S <= D(0) WHEN 0,
     D(1) WHEN 1,
     D(2) WHEN 2,
     D(3) WHEN 3;
END CIR;