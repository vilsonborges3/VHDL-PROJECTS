ENTITY LATCHRS IS 
PORT (SETA, RESETA : IN BIT;
		Q: BUFFER BIT);
END LATCHRS;

ARCHITECTURE CIR OF LATCHRS IS
BEGIN 

	PROCESS (SETA, RESETA)
	BEGIN
		IF SETA = '1' THEN Q <= '1';
		ELSIF RESETA = '1' THEN Q <= '0';
		ELSE Q <= Q;
		END IF;
	END PROCESS;
END CIR; 