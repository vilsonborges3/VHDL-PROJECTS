--PROVA 2 VILSON BORGES - 12011EAU020

ENTITY CIRCUITO IS 
PORT ( CLOCK, INICIA : IN BIT;
       MAIOR, IGUAL, MENOR: OUT BIT);
END CIRCUITO;

ARCHITECTURE CIR1 OF CIRCUITO IS

COMPONENT FLIPFLOP
PORT ( PRN, CLRN, CLKN, J, K : IN BIT ;
       Q : BUFFER BIT ) ;
END COMPONENT ;

SIGNAL Q0, Q1, Q2, Q3, Q4, Q5: BIT;
SIGNAL A0, A1: BIT;
SIGNAL AUX1: BIT;
SIGNAL AUX2, AUX3: BIT_VECTOR (3 DOWNTO 0);

BEGIN
--PROJETO FLIP-FLPS
FF0 : FLIPFLOP PORT MAP (PRN => INICIA, CLRN => '1', CLKN => CLOCK, J => Q0 AND (NOT Q1),  K => '1',Q => Q2) ;
FF1 : FLIPFLOP PORT MAP (PRN => INICIA, CLRN => '1', CLKN => CLOCK, J => '1',   K => '1',     Q => Q1) ;
FF2 : FLIPFLOP PORT MAP (PRN => INICIA, CLRN => '1', CLKN => CLOCK, J => '1',  K => Q2,     Q => Q0) ;

AUX1 <= (NOT((NOT Q3 ) AND Q4 AND Q5)) AND INICIA;

FF3 : FLIPFLOP PORT MAP (PRN => AUX1, CLRN => '1', CLKN => CLOCK,  J => '1', K => '1', Q => Q3);
FF4 : FLIPFLOP PORT MAP (PRN => '1', CLRN => AUX1, CLKN => Q3,  J => '1',K => '1', Q => Q4);
FF5 : FLIPFLOP PORT MAP (PRN => '1', CLRN => AUX1, CLKN => Q4,  J => '1',K => '1', Q => Q5);

--PROJETO DO CIRCUITO 1
AUX2 <= Q2&Q1&Q0&Q3;
WITH AUX2 SELECT
A1 <= '1' WHEN "0000",
	 '0' WHEN "0001",
	 '1' WHEN "0010",
	 '1' WHEN "0011",
	 '0' WHEN "0100",
	 '1' WHEN "0101",
	 '1' WHEN "0110",
	 '1' WHEN "0111",
	 '1' WHEN "1000",
	 '1' WHEN "1001",
	 '1' WHEN "1010",
	 '0' WHEN "1011",
	 '0' WHEN "1100",
	 '0' WHEN "1101",
	 '1' WHEN "1110",
	 '1' WHEN "1111";
	 
WITH AUX2 SELECT
A0 <= '0' WHEN "0000",
	 '1' WHEN "0001",
	 '0' WHEN "0010",
	 '0' WHEN "0011",
	 '1' WHEN "0100",
	 '0' WHEN "0101",
	 '1' WHEN "0110",
	 '0' WHEN "0111",
	 '1' WHEN "1000",
	 '0' WHEN "1001",
	 '1' WHEN "1010",
	 '1' WHEN "1011",
	 '0' WHEN "1100",
	 '1' WHEN "1101",
	 '1' WHEN "1110",
	 '0' WHEN "1111";

--PROJETO DO CIRCUITO COMPARADOR 
AUX3 <= A1&A0&Q4&Q5;
WITH AUX3 SELECT
MAIOR <= '0' WHEN "0000",
		 '0' WHEN "0001",
		 '0' WHEN "0010",
		 '0' WHEN "0011",
		 '1' WHEN "0100",
		 '0' WHEN "0101",
		 '0' WHEN "0110",
		 '0' WHEN "0111",
		 '1' WHEN "1000",
		 '1' WHEN "1001",
		 '0' WHEN "1010",
		 '0' WHEN "1011",
		 '1' WHEN "1100",
		 '1' WHEN "1101",
		 '1' WHEN "1110",
		 '0' WHEN "1111";

WITH AUX3 SELECT
IGUAL <= '1' WHEN "0000",
		 '0' WHEN "0001",
		 '0' WHEN "0010",
		 '0' WHEN "0011",
		 '0' WHEN "0100",
		 '1' WHEN "0101",
		 '0' WHEN "0110",
		 '0' WHEN "0111",
		 '0' WHEN "1000",
		 '0' WHEN "1001",
		 '1' WHEN "1010",
		 '0' WHEN "1011",
		 '0' WHEN "1100",
		 '0' WHEN "1101",
		 '0' WHEN "1110",
		 '1' WHEN "1111";
		 
WITH AUX3 SELECT
MENOR <= '0' WHEN "0000",
		 '1' WHEN "0001",
		 '1' WHEN "0010",
		 '1' WHEN "0011",
		 '0' WHEN "0100",
		 '0' WHEN "0101",
		 '1' WHEN "0110",
		 '1' WHEN "0111",
		 '0' WHEN "1000",
		 '0' WHEN "1001",
		 '0' WHEN "1010",
		 '1' WHEN "1011",
		 '0' WHEN "1100",
		 '0' WHEN "1101",
		 '0' WHEN "1110",
		 '0' WHEN "1111";
END CIR1;



-- PROJETO DO FLIP FLOP JK MESTRE-ESCRAVO COM PRESET E CLEAR.

ENTITY FLIPFLOP IS
PORT ( PRN, CLRN, CLKN, J, K : IN BIT ;
       Q : BUFFER BIT ) ;
END FLIPFLOP ;

ARCHITECTURE CIR OF FLIPFLOP IS
BEGIN
	PROCESS ( PRN, CLRN, CLKN )
	BEGIN
		IF     PRN = '0' THEN Q <= '1' ;
		ELSIF CLRN = '0' THEN Q <= '0' ;
		ELSIF CLKN = '0' AND CLKN 'EVENT THEN 
			IF    J = '1' AND K = '1' THEN Q <= NOT Q ;
			ELSIF J = '1' AND K = '0' THEN Q <= '1' ;
			ELSIF J = '0' AND K = '1' THEN Q <= '0' ;
            END IF;
        END IF ;
    END PROCESS ;
    Q <= Q ;

END CIR ;