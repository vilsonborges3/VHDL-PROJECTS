
ENTITY M12011EAU020 IS
PORT (D0, D1, D2, D3 : IN BIT ;
		A0, A1 : IN BIT;
		B0, B1, B2: IN BIT;
		S0, S1, S2, S3, S4, S5, S6, S7: OUT BIT );
END M12011EAU020 ;

ARCHITECTURE CIR OF M12011EAU020 IS 

SIGNAL E : BIT;
SIGNAL AA : BIT_VECTOR (1 DOWNTO 0) ;
SIGNAL BB : BIT_VECTOR (2 DOWNTO 0) ;


BEGIN 
AA <= A1 & A0; 
BB <= B2 & B1 & B0;
WITH AA SELECT

E <= D0 WHEN "00",
     D1 WHEN "01",
     D2 WHEN "10",
     D3 WHEN "11";

S0 <= E WHEN BB = "000" ELSE '1';
S1 <= E WHEN BB = "001" ELSE '1';
S2 <= E WHEN BB = "010" ELSE '1';
S3 <= E WHEN BB = "011" ELSE '1';
S4 <= E WHEN BB = "100" ELSE '1';
S5 <= E WHEN BB = "101" ELSE '1';
S6 <= E WHEN BB = "110" ELSE '1';
S7 <= E WHEN BB = "111" ELSE '1';
END CIR;