-- TRABALHO 08
-- VILSON B 12011EAU020

ENTITY CIRCUITO IS
PORT ( INICIA, CLOCK : IN BIT ;
       S : OUT BIT ) ;
END CIRCUITO ;

ARCHITECTURE CIR1 OF CIRCUITO IS

COMPONENT FLIPFLOP
PORT ( PRN, CLRN, CLKN, J, K : IN BIT ;
       Q : BUFFER BIT ) ;
END COMPONENT ;

SIGNAL S1, S2: BIT;
SIGNAL AUX1, AUX2, AUX3, AUX4: BIT;
SIGNAL Q0, Q1, Q2, Q3, Q4, Q5: BIT;
SIGNAL A : BIT_VECTOR ( 2 DOWNTO 0);
BEGIN

WITH A SELECT
   S1<='0' WHEN "000",
	   '1' WHEN "001",
	   '0' WHEN "010",
	   '1' WHEN "011",
	   '0' WHEN "100",
	   '1' WHEN "101",
	   '1' WHEN "110",
	   '1' WHEN "111";

A(0)<=Q0;
A(1)<=Q1;
A(2)<=Q3;

AUX1 <= NOT(NOT(Q2) AND Q0 AND NOT(Q1)) AND INICIA;
AUX2 <= Q4 XOR Q3;


FF0 : FLIPFLOP PORT MAP (PRN => '1', CLRN => AUX1, CLKN => CLOCK, J => '1',  K => '1',     Q => Q0) ;
FF1 : FLIPFLOP PORT MAP (PRN => AUX1, CLRN => '1' , CLKN => NOT(Q0), J => '1',  K => '1',     Q => Q1) ;
FF2 : FLIPFLOP PORT MAP (PRN => AUX1, CLRN => '1' , CLKN => NOT(Q1), J => '1',  K => '1',     Q => Q2) ;

FF3 : FLIPFLOP PORT MAP (PRN => '1', CLRN => INICIA , CLKN => AUX1, J => '1',  K => '1',     Q => Q3) ;
FF4 : FLIPFLOP PORT MAP (PRN => '1', CLRN => INICIA , CLKN => AUX1, J => Q3,  K => Q3,     Q => Q4) ;
FF5 : FLIPFLOP PORT MAP (PRN => '1', CLRN => INICIA , CLKN => AUX1, J => AUX2,  K => AUX2,     Q => Q5) ;

AUX3 <= Q4 XNOR Q5;
AUX4 <= NOT (S1 OR S2);
S <= NOT (AUX4 AND AUX3);

END CIR1 ;

-- PROJETO DO FLIP FLOP JK MESTRE-ESCRAVO COM PRESET E CLEAR.

ENTITY FLIPFLOP IS
PORT ( PRN, CLRN, CLKN, J, K : IN BIT ;
       Q : BUFFER BIT ) ;
END FLIPFLOP ;

ARCHITECTURE CIR OF FLIPFLOP IS
BEGIN
	PROCESS ( PRN, CLRN, CLKN )
	BEGIN
		IF     PRN = '0' THEN Q <= '1' ;
		ELSIF CLRN = '0' THEN Q <= '0' ;
		ELSIF CLKN = '0' AND CLKN 'EVENT THEN 
			IF    J = '1' AND K = '1' THEN Q <= NOT Q ;
			ELSIF J = '1' AND K = '0' THEN Q <= '1' ;
			ELSIF J = '0' AND K = '1' THEN Q <= '0' ;
            END IF;
        END IF ;
    END PROCESS ;
    Q <= Q ;

END CIR ;